module IF_Stage_Reg (
  input clk, rst, freeze, flush, 
  input[31:0] PCIn, Instrution_in, 
  output reg[31:0] PC, Instruction
  );
  always @ (posedge clk) begin
    if (rst) begin
      {PC} <= 0;
      {Instruction} <= 32'b0;
    end
    else begin
      PC <= PCIn;
      {Instruction} <= Instruction_in;
    end
  end
endmodule